interface ubus_s_if;

	logic ubus_clock;
	logic ubus_reset;
	logic [15:0] ubus_addr;
	logic [2:0] ubus_size;
	logic ubus_read;
	logic ubus_write;
	logic ubus_bip;
	logic [7:0] ubus_data;
	logic ubus_wait;
	logic ubus_error;




endinterface
